module sad (input wire [64-1:0] crt_frame,
                  input wire [64-1:0] pre_frame,
                  output wire [14+4-1:0] sad,
                  );
    
endmodule
