module core_ctrl (
    
);
    
endmodule