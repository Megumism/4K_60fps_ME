module sad (
    input wire clk,
    input wire rst,
    input wire crt_keep,
    input wire [64-1:0] crt_frame,
                  input wire [64-1:0] pre_frame,
                  output wire [14-1:0] sad
                //   output wire [4-1:0] motion_vec_y
                  );
    
endmodule
