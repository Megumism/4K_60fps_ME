module sad (input wire clk,
            input wire rst_n,
            input wire crt_keep,
            input wire [64-1:0] pre_frame,
            input wire [64-1:0] crt_frame,
            output reg [14-1:0] sad_data);
    
    wire [8-1:0] crt_pixel_o_00, pre_pixel_o_00, ad_00;
    pe pe_00(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep) 
       ,.crt_pixel_i(crt_frame[63:56])
       ,.pre_pixel_i(pre_frame[63:56])
       ,.crt_pixel_o(crt_pixel_o_00)
       ,.pre_pixel_o(pre_pixel_o_00)
       ,.ad(ad_00)
    );

    wire [8-1:0] crt_pixel_o_01, pre_pixel_o_01, ad_01;
    pe pe_01(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep) 
       ,.crt_pixel_i(crt_frame[55:48])
       ,.pre_pixel_i(pre_frame[55:48])
       ,.crt_pixel_o(crt_pixel_o_01)
       ,.pre_pixel_o(pre_pixel_o_01)
       ,.ad(ad_01)
       
    );

    wire [8-1:0] crt_pixel_o_02, pre_pixel_o_02, ad_02;
    pe pe_02(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep) 
       ,.crt_pixel_i(crt_frame[47:40])
       ,.pre_pixel_i(pre_frame[47:40])
       ,.crt_pixel_o(crt_pixel_o_02)
       ,.pre_pixel_o(pre_pixel_o_02)
       ,.ad(ad_02)
       
    );

    wire [8-1:0] crt_pixel_o_03, pre_pixel_o_03, ad_03;
    pe pe_03(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep) 
       ,.crt_pixel_i(crt_frame[39:32])
       ,.pre_pixel_i(pre_frame[39:32])
       ,.crt_pixel_o(crt_pixel_o_03)
       ,.pre_pixel_o(pre_pixel_o_03)
       ,.ad(ad_03)
       
    );

    wire [8-1:0] crt_pixel_o_04, pre_pixel_o_04, ad_04;
    pe pe_04(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep) 
       ,.crt_pixel_i(crt_frame[31:24])
       ,.pre_pixel_i(pre_frame[31:24])
       ,.crt_pixel_o(crt_pixel_o_04)
       ,.pre_pixel_o(pre_pixel_o_04)
       ,.ad(ad_04)
       
    );

    wire [8-1:0] crt_pixel_o_05, pre_pixel_o_05, ad_05;
    pe pe_05(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep) 
       ,.crt_pixel_i(crt_frame[23:16])
       ,.pre_pixel_i(pre_frame[23:16])
       ,.crt_pixel_o(crt_pixel_o_05)
       ,.pre_pixel_o(pre_pixel_o_05)
       ,.ad(ad_05)
       
    );

    wire [8-1:0] crt_pixel_o_06, pre_pixel_o_06, ad_06;
    pe pe_06(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep) 
       ,.crt_pixel_i(crt_frame[15:8])
       ,.pre_pixel_i(pre_frame[15:8])
       ,.crt_pixel_o(crt_pixel_o_06)
       ,.pre_pixel_o(pre_pixel_o_06)
       ,.ad(ad_06)
       
    );

    wire [8-1:0] crt_pixel_o_07, pre_pixel_o_07, ad_07;
    pe pe_07(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep) 
       ,.crt_pixel_i(crt_frame[7:0])
       ,.pre_pixel_i(pre_frame[7:0])
       ,.crt_pixel_o(crt_pixel_o_07)
       ,.pre_pixel_o(pre_pixel_o_07)
       ,.ad(ad_07)
       
    );

    wire [8-1:0] crt_pixel_o_10, pre_pixel_o_10, ad_10;
    pe pe_10(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep) 
       ,.crt_pixel_i(crt_pixel_o_00)
       ,.pre_pixel_i(pre_pixel_o_00)
       ,.crt_pixel_o(crt_pixel_o_10)
       ,.pre_pixel_o(pre_pixel_o_10)
       ,.ad(ad_10)
       
    );

    wire [8-1:0] crt_pixel_o_11, pre_pixel_o_11, ad_11;
    pe pe_11(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep) 
       ,.crt_pixel_i(crt_pixel_o_01)
       ,.pre_pixel_i(pre_pixel_o_01)
       ,.crt_pixel_o(crt_pixel_o_11)
       ,.pre_pixel_o(pre_pixel_o_11)
       ,.ad(ad_11)
       
    );

    wire [8-1:0] crt_pixel_o_12, pre_pixel_o_12, ad_12;
    pe pe_12(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep) 
       ,.crt_pixel_i(crt_pixel_o_02)
       ,.pre_pixel_i(pre_pixel_o_02)
       ,.crt_pixel_o(crt_pixel_o_12)
       ,.pre_pixel_o(pre_pixel_o_12)
       ,.ad(ad_12)
       
    );

    wire [8-1:0] crt_pixel_o_13, pre_pixel_o_13, ad_13;
    pe pe_13(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep)
       ,.crt_pixel_i(crt_pixel_o_03)
       ,.pre_pixel_i(pre_pixel_o_03)
       ,.crt_pixel_o(crt_pixel_o_13)
       ,.pre_pixel_o(pre_pixel_o_13)
       ,.ad(ad_13)
       
    );

    wire [8-1:0] crt_pixel_o_14, pre_pixel_o_14, ad_14;
    pe pe_14(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep) 
       ,.crt_pixel_i(crt_pixel_o_04)
       ,.pre_pixel_i(pre_pixel_o_04)
       ,.crt_pixel_o(crt_pixel_o_14)
       ,.pre_pixel_o(pre_pixel_o_14)
       ,.ad(ad_14)
       
    );

    wire [8-1:0] crt_pixel_o_15, pre_pixel_o_15, ad_15;
    pe pe_15(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep) 
       ,.crt_pixel_i(crt_pixel_o_05)
       ,.pre_pixel_i(pre_pixel_o_05)
       ,.crt_pixel_o(crt_pixel_o_15)
       ,.pre_pixel_o(pre_pixel_o_15)
       ,.ad(ad_15)
       
    );

    wire [8-1:0] crt_pixel_o_16, pre_pixel_o_16, ad_16;
    pe pe_16(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep) 
       ,.crt_pixel_i(crt_pixel_o_06)
       ,.pre_pixel_i(pre_pixel_o_06)
       ,.crt_pixel_o(crt_pixel_o_16)
       ,.pre_pixel_o(pre_pixel_o_16)
       ,.ad(ad_16)
       
    );

    wire [8-1:0] crt_pixel_o_17, pre_pixel_o_17, ad_17;
    pe pe_17(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep) 
       ,.crt_pixel_i(crt_pixel_o_07)
       ,.pre_pixel_i(pre_pixel_o_07)
       ,.crt_pixel_o(crt_pixel_o_17)
       ,.pre_pixel_o(pre_pixel_o_17)
       ,.ad(ad_17)
       
    );

    wire [8-1:0] crt_pixel_o_20, pre_pixel_o_20, ad_20;
    pe pe_20(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep) 
       ,.crt_pixel_i(crt_pixel_o_10)
       ,.pre_pixel_i(pre_pixel_o_10)
       ,.crt_pixel_o(crt_pixel_o_20)
       ,.pre_pixel_o(pre_pixel_o_20)
       ,.ad(ad_20)
       
    );

    wire [8-1:0] crt_pixel_o_21, pre_pixel_o_21, ad_21;
    pe pe_21(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep) 
       ,.crt_pixel_i(crt_pixel_o_11)
       ,.pre_pixel_i(pre_pixel_o_11)
       ,.crt_pixel_o(crt_pixel_o_21)
       ,.pre_pixel_o(pre_pixel_o_21)
       ,.ad(ad_21)
       
    );

    wire [8-1:0] crt_pixel_o_22, pre_pixel_o_22, ad_22;
    pe pe_22(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep) 
       ,.crt_pixel_i(crt_pixel_o_12)
       ,.pre_pixel_i(pre_pixel_o_12)
       ,.crt_pixel_o(crt_pixel_o_22)
       ,.pre_pixel_o(pre_pixel_o_22)
       ,.ad(ad_22)
       
    );

    wire [8-1:0] crt_pixel_o_23, pre_pixel_o_23, ad_23;
    pe pe_23(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep) 
       ,.crt_pixel_i(crt_pixel_o_13)
       ,.pre_pixel_i(pre_pixel_o_13)
       ,.crt_pixel_o(crt_pixel_o_23)
       ,.pre_pixel_o(pre_pixel_o_23)
       ,.ad(ad_23)
       
    );

    wire [8-1:0] crt_pixel_o_24, pre_pixel_o_24, ad_24;
    pe pe_24(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep) 
       ,.crt_pixel_i(crt_pixel_o_14)
       ,.pre_pixel_i(pre_pixel_o_14)
       ,.crt_pixel_o(crt_pixel_o_24)
       ,.pre_pixel_o(pre_pixel_o_24)
       ,.ad(ad_24)
       
    );

    wire [8-1:0] crt_pixel_o_25, pre_pixel_o_25, ad_25;
    pe pe_25(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep) 
       ,.crt_pixel_i(crt_pixel_o_15)
       ,.pre_pixel_i(pre_pixel_o_15)
       ,.crt_pixel_o(crt_pixel_o_25)
       ,.pre_pixel_o(pre_pixel_o_25)
       ,.ad(ad_25)
       
    );

    wire [8-1:0] crt_pixel_o_26, pre_pixel_o_26, ad_26;
    pe pe_26(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep) 
       ,.crt_pixel_i(crt_pixel_o_16)
       ,.pre_pixel_i(pre_pixel_o_16)
       ,.crt_pixel_o(crt_pixel_o_26)
       ,.pre_pixel_o(pre_pixel_o_26)
       ,.ad(ad_26)
       
    );

    wire [8-1:0] crt_pixel_o_27, pre_pixel_o_27, ad_27;
    pe pe_27(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep) 
       ,.crt_pixel_i(crt_pixel_o_17)
       ,.pre_pixel_i(pre_pixel_o_17)
       ,.crt_pixel_o(crt_pixel_o_27)
       ,.pre_pixel_o(pre_pixel_o_27)
       ,.ad(ad_27)
       
    );

    wire [8-1:0] crt_pixel_o_30, pre_pixel_o_30, ad_30;
    pe pe_30(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep) 
       ,.crt_pixel_i(crt_pixel_o_20)
       ,.pre_pixel_i(pre_pixel_o_20)
       ,.crt_pixel_o(crt_pixel_o_30)
       ,.pre_pixel_o(pre_pixel_o_30)
       ,.ad(ad_30)
       
    );

    wire [8-1:0] crt_pixel_o_31, pre_pixel_o_31, ad_31;
    pe pe_31(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep) 
       ,.crt_pixel_i(crt_pixel_o_21)
       ,.pre_pixel_i(pre_pixel_o_21)
       ,.crt_pixel_o(crt_pixel_o_31)
       ,.pre_pixel_o(pre_pixel_o_31)
       ,.ad(ad_31)
       
    );

    wire [8-1:0] crt_pixel_o_32, pre_pixel_o_32, ad_32;
    pe pe_32(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep) 
       ,.crt_pixel_i(crt_pixel_o_22)
       ,.pre_pixel_i(pre_pixel_o_22)
       ,.crt_pixel_o(crt_pixel_o_32)
       ,.pre_pixel_o(pre_pixel_o_32)
       ,.ad(ad_32)
       
    );

    wire [8-1:0] crt_pixel_o_33, pre_pixel_o_33, ad_33;
    pe pe_33(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep)
       ,.crt_pixel_i(crt_pixel_o_23)
       ,.pre_pixel_i(pre_pixel_o_23)
       ,.crt_pixel_o(crt_pixel_o_33)
       ,.pre_pixel_o(pre_pixel_o_33)
       ,.ad(ad_33)
       
    );

    wire [8-1:0] crt_pixel_o_34, pre_pixel_o_34, ad_34;
    pe pe_34(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep) 
       ,.crt_pixel_i(crt_pixel_o_24)
       ,.pre_pixel_i(pre_pixel_o_24)
       ,.crt_pixel_o(crt_pixel_o_34)
       ,.pre_pixel_o(pre_pixel_o_34)
       ,.ad(ad_34)
       
    );

    wire [8-1:0] crt_pixel_o_35, pre_pixel_o_35, ad_35;
    pe pe_35(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep) 
       ,.crt_pixel_i(crt_pixel_o_25)
       ,.pre_pixel_i(pre_pixel_o_25)
       ,.crt_pixel_o(crt_pixel_o_35)
       ,.pre_pixel_o(pre_pixel_o_35)
       ,.ad(ad_35)
       
    );

    wire [8-1:0] crt_pixel_o_36, pre_pixel_o_36, ad_36;
    pe pe_36(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep) 
       ,.crt_pixel_i(crt_pixel_o_26)
       ,.pre_pixel_i(pre_pixel_o_26)
       ,.crt_pixel_o(crt_pixel_o_36)
       ,.pre_pixel_o(pre_pixel_o_36)
       ,.ad(ad_36)
       
    );

    wire [8-1:0] crt_pixel_o_37, pre_pixel_o_37, ad_37;
    pe pe_37(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep) 
       ,.crt_pixel_i(crt_pixel_o_27)
       ,.pre_pixel_i(pre_pixel_o_27)
       ,.crt_pixel_o(crt_pixel_o_37)
       ,.pre_pixel_o(pre_pixel_o_37)
       ,.ad(ad_37)
       
    );

    wire [8-1:0] crt_pixel_o_40, pre_pixel_o_40, ad_40;
    pe pe_40(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep) 
       ,.crt_pixel_i(crt_pixel_o_30)
       ,.pre_pixel_i(pre_pixel_o_30)
       ,.crt_pixel_o(crt_pixel_o_40)
       ,.pre_pixel_o(pre_pixel_o_40)
       ,.ad(ad_40)
       
    );

    wire [8-1:0] crt_pixel_o_41, pre_pixel_o_41, ad_41;
    pe pe_41(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep) 
       ,.crt_pixel_i(crt_pixel_o_31)
       ,.pre_pixel_i(pre_pixel_o_31)
       ,.crt_pixel_o(crt_pixel_o_41)
       ,.pre_pixel_o(pre_pixel_o_41)
       ,.ad(ad_41)
       
    );

    wire [8-1:0] crt_pixel_o_42, pre_pixel_o_42, ad_42;
    pe pe_42(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep) 
       ,.crt_pixel_i(crt_pixel_o_32)
       ,.pre_pixel_i(pre_pixel_o_32)
       ,.crt_pixel_o(crt_pixel_o_42)
       ,.pre_pixel_o(pre_pixel_o_42)
       ,.ad(ad_42)
       
    );

    wire [8-1:0] crt_pixel_o_43, pre_pixel_o_43, ad_43;
    pe pe_43(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep)
       ,.crt_pixel_i(crt_pixel_o_33)
       ,.pre_pixel_i(pre_pixel_o_33)
       ,.crt_pixel_o(crt_pixel_o_43)
       ,.pre_pixel_o(pre_pixel_o_43)
       ,.ad(ad_43)
       
    );

    wire [8-1:0] crt_pixel_o_44, pre_pixel_o_44, ad_44;
    pe pe_44(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep) 
       ,.crt_pixel_i(crt_pixel_o_34)
       ,.pre_pixel_i(pre_pixel_o_34)
       ,.crt_pixel_o(crt_pixel_o_44)
       ,.pre_pixel_o(pre_pixel_o_44)
       ,.ad(ad_44)
       
    );

    wire [8-1:0] crt_pixel_o_45, pre_pixel_o_45, ad_45;
    pe pe_45(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep) 
       ,.crt_pixel_i(crt_pixel_o_35)
       ,.pre_pixel_i(pre_pixel_o_35)
       ,.crt_pixel_o(crt_pixel_o_45)
       ,.pre_pixel_o(pre_pixel_o_45)
       ,.ad(ad_45)
       
    );

    wire [8-1:0] crt_pixel_o_46, pre_pixel_o_46, ad_46;
    pe pe_46(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep) 
       ,.crt_pixel_i(crt_pixel_o_36)
       ,.pre_pixel_i(pre_pixel_o_36)
       ,.crt_pixel_o(crt_pixel_o_46)
       ,.pre_pixel_o(pre_pixel_o_46)
       ,.ad(ad_46)
       
    );

    wire [8-1:0] crt_pixel_o_47, pre_pixel_o_47, ad_47;
    pe pe_47(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep) 
       ,.crt_pixel_i(crt_pixel_o_37)
       ,.pre_pixel_i(pre_pixel_o_37)
       ,.crt_pixel_o(crt_pixel_o_47)
       ,.pre_pixel_o(pre_pixel_o_47)
       ,.ad(ad_47)
       
    );

    wire [8-1:0] crt_pixel_o_50, pre_pixel_o_50, ad_50;
    pe pe_50(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep) 
       ,.crt_pixel_i(crt_pixel_o_40)
       ,.pre_pixel_i(pre_pixel_o_40)
       ,.crt_pixel_o(crt_pixel_o_50)
       ,.pre_pixel_o(pre_pixel_o_50)
       ,.ad(ad_50)
       
    );

    wire [8-1:0] crt_pixel_o_51, pre_pixel_o_51, ad_51;
    pe pe_51(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep) 
       ,.crt_pixel_i(crt_pixel_o_41)
       ,.pre_pixel_i(pre_pixel_o_41)
       ,.crt_pixel_o(crt_pixel_o_51)
       ,.pre_pixel_o(pre_pixel_o_51)
       ,.ad(ad_51)
       
    );

    wire [8-1:0] crt_pixel_o_52, pre_pixel_o_52, ad_52;
    pe pe_52(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep) 
       ,.crt_pixel_i(crt_pixel_o_42)
       ,.pre_pixel_i(pre_pixel_o_42)
       ,.crt_pixel_o(crt_pixel_o_52)
       ,.pre_pixel_o(pre_pixel_o_52)
       ,.ad(ad_52)
       
    );

    wire [8-1:0] crt_pixel_o_53, pre_pixel_o_53, ad_53;
    pe pe_53(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep)
       ,.crt_pixel_i(crt_pixel_o_43)
       ,.pre_pixel_i(pre_pixel_o_43)
       ,.crt_pixel_o(crt_pixel_o_53)
       ,.pre_pixel_o(pre_pixel_o_53)
       ,.ad(ad_53)
       
    );

    wire [8-1:0] crt_pixel_o_54, pre_pixel_o_54, ad_54;
    pe pe_54(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep) 
       ,.crt_pixel_i(crt_pixel_o_44)
       ,.pre_pixel_i(pre_pixel_o_44)
       ,.crt_pixel_o(crt_pixel_o_54)
       ,.pre_pixel_o(pre_pixel_o_54)
       ,.ad(ad_54)
       
    );

    wire [8-1:0] crt_pixel_o_55, pre_pixel_o_55, ad_55;
    pe pe_55(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep) 
       ,.crt_pixel_i(crt_pixel_o_45)
       ,.pre_pixel_i(pre_pixel_o_45)
       ,.crt_pixel_o(crt_pixel_o_55)
       ,.pre_pixel_o(pre_pixel_o_55)
       ,.ad(ad_55)
       
    );

    wire [8-1:0] crt_pixel_o_56, pre_pixel_o_56, ad_56;
    pe pe_56(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep) 
       ,.crt_pixel_i(crt_pixel_o_46)
       ,.pre_pixel_i(pre_pixel_o_46)
       ,.crt_pixel_o(crt_pixel_o_56)
       ,.pre_pixel_o(pre_pixel_o_56)
       ,.ad(ad_56)
       
    );

    wire [8-1:0] crt_pixel_o_57, pre_pixel_o_57, ad_57;
    pe pe_57(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep) 
       ,.crt_pixel_i(crt_pixel_o_47)
       ,.pre_pixel_i(pre_pixel_o_47)
       ,.crt_pixel_o(crt_pixel_o_57)
       ,.pre_pixel_o(pre_pixel_o_57)
       ,.ad(ad_57)
       
    );

    wire [8-1:0] crt_pixel_o_60, pre_pixel_o_60, ad_60;
    pe pe_60(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep) 
       ,.crt_pixel_i(crt_pixel_o_50)
       ,.pre_pixel_i(pre_pixel_o_50)
       ,.crt_pixel_o(crt_pixel_o_60)
       ,.pre_pixel_o(pre_pixel_o_60)
       ,.ad(ad_60)
       
    );

    wire [8-1:0] crt_pixel_o_61, pre_pixel_o_61, ad_61;
    pe pe_61(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep) 
       ,.crt_pixel_i(crt_pixel_o_51)
       ,.pre_pixel_i(pre_pixel_o_51)
       ,.crt_pixel_o(crt_pixel_o_61)
       ,.pre_pixel_o(pre_pixel_o_61)
       ,.ad(ad_61)
       
    );

    wire [8-1:0] crt_pixel_o_62, pre_pixel_o_62, ad_62;
    pe pe_62(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep) 
       ,.crt_pixel_i(crt_pixel_o_52)
       ,.pre_pixel_i(pre_pixel_o_52)
       ,.crt_pixel_o(crt_pixel_o_62)
       ,.pre_pixel_o(pre_pixel_o_62)
       ,.ad(ad_62)
       
    );

    wire [8-1:0] crt_pixel_o_63, pre_pixel_o_63, ad_63;
    pe pe_63(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep) 
       ,.crt_pixel_i(crt_pixel_o_53)
       ,.pre_pixel_i(pre_pixel_o_53)
       ,.crt_pixel_o(crt_pixel_o_63)
       ,.pre_pixel_o(pre_pixel_o_63)
       ,.ad(ad_63)
       
    );

    wire [8-1:0] crt_pixel_o_64, pre_pixel_o_64, ad_64;
    pe pe_64(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep) 
       ,.crt_pixel_i(crt_pixel_o_54)
       ,.pre_pixel_i(pre_pixel_o_54)
       ,.crt_pixel_o(crt_pixel_o_64)
       ,.pre_pixel_o(pre_pixel_o_64)
       ,.ad(ad_64)
       
    );

    wire [8-1:0] crt_pixel_o_65, pre_pixel_o_65, ad_65;
    pe pe_65(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep) 
       ,.crt_pixel_i(crt_pixel_o_55)
       ,.pre_pixel_i(pre_pixel_o_55)
       ,.crt_pixel_o(crt_pixel_o_65)
       ,.pre_pixel_o(pre_pixel_o_65)
       ,.ad(ad_65)
       
    );

    wire [8-1:0] crt_pixel_o_66, pre_pixel_o_66, ad_66;
    pe pe_66(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep) 
       ,.crt_pixel_i(crt_pixel_o_56)
       ,.pre_pixel_i(pre_pixel_o_56)
       ,.crt_pixel_o(crt_pixel_o_66)
       ,.pre_pixel_o(pre_pixel_o_66)
       ,.ad(ad_66)
       
    );

    wire [8-1:0] crt_pixel_o_67, pre_pixel_o_67, ad_67;
    pe pe_67(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep) 
       ,.crt_pixel_i(crt_pixel_o_57)
       ,.pre_pixel_i(pre_pixel_o_57)
       ,.crt_pixel_o(crt_pixel_o_67)
       ,.pre_pixel_o(pre_pixel_o_67)
       ,.ad(ad_67)
       
    );

    wire [8-1:0] crt_pixel_o_70, pre_pixel_o_70, ad_70;
    pe pe_70(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep) 
       ,.crt_pixel_i(crt_pixel_o_60)
       ,.pre_pixel_i(pre_pixel_o_60)
       ,.crt_pixel_o(crt_pixel_o_70)
       ,.pre_pixel_o(pre_pixel_o_70)
       ,.ad(ad_70)
       
    );

    wire [8-1:0] crt_pixel_o_71, pre_pixel_o_71, ad_71;
    pe pe_71(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep) 
       ,.crt_pixel_i(crt_pixel_o_61)
       ,.pre_pixel_i(pre_pixel_o_61)
       ,.crt_pixel_o(crt_pixel_o_71)
       ,.pre_pixel_o(pre_pixel_o_71)
       ,.ad(ad_71)
       
    );

    wire [8-1:0] crt_pixel_o_72, pre_pixel_o_72, ad_72;
    pe pe_72(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep) 
       ,.crt_pixel_i(crt_pixel_o_62)
       ,.pre_pixel_i(pre_pixel_o_62)
       ,.crt_pixel_o(crt_pixel_o_72)
       ,.pre_pixel_o(pre_pixel_o_72)
       ,.ad(ad_72)
       
    );

    wire [8-1:0] crt_pixel_o_73, pre_pixel_o_73, ad_73;
    pe pe_73(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep) 
       ,.crt_pixel_i(crt_pixel_o_63)
       ,.pre_pixel_i(pre_pixel_o_63)
       ,.crt_pixel_o(crt_pixel_o_73)
       ,.pre_pixel_o(pre_pixel_o_73)
       ,.ad(ad_73)
       
    );

    wire [8-1:0] crt_pixel_o_74, pre_pixel_o_74, ad_74;
    pe pe_74(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep) 
       ,.crt_pixel_i(crt_pixel_o_64)
       ,.pre_pixel_i(pre_pixel_o_64)
       ,.crt_pixel_o(crt_pixel_o_74)
       ,.pre_pixel_o(pre_pixel_o_74)
       ,.ad(ad_74)
       
    );

    wire [8-1:0] crt_pixel_o_75, pre_pixel_o_75, ad_75;
    pe pe_75(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep) 
       ,.crt_pixel_i(crt_pixel_o_65)
       ,.pre_pixel_i(pre_pixel_o_65)
       ,.crt_pixel_o(crt_pixel_o_75)
       ,.pre_pixel_o(pre_pixel_o_75)
       ,.ad(ad_75)
       
    );

    wire [8-1:0] crt_pixel_o_76, pre_pixel_o_76, ad_76;
    pe pe_76(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep) 
       ,.crt_pixel_i(crt_pixel_o_66)
       ,.pre_pixel_i(pre_pixel_o_66)
       ,.crt_pixel_o(crt_pixel_o_76)
       ,.pre_pixel_o(pre_pixel_o_76)
       ,.ad(ad_76)
       
    );

    wire [8-1:0] crt_pixel_o_77, pre_pixel_o_77, ad_77;
    pe pe_77(
        .clk(clk)
       ,.rst_n(rst_n)
       ,.crt_keep(crt_keep) 
       ,.crt_pixel_i(crt_pixel_o_67)
       ,.pre_pixel_i(pre_pixel_o_67)
       ,.crt_pixel_o(crt_pixel_o_77)
       ,.pre_pixel_o(pre_pixel_o_77)
       ,.ad(ad_77)
       
    );

    //adder_tree
    wire [9-1:0] add_0_00;
    wire [9-1:0] add_0_01;
    wire [9-1:0] add_0_02;
    wire [9-1:0] add_0_03;
    wire [9-1:0] add_0_04;
    wire [9-1:0] add_0_05;
    wire [9-1:0] add_0_06;
    wire [9-1:0] add_0_07;
    wire [9-1:0] add_0_08;
    wire [9-1:0] add_0_09;
    wire [9-1:0] add_0_10;
    wire [9-1:0] add_0_11;
    wire [9-1:0] add_0_12;
    wire [9-1:0] add_0_13;
    wire [9-1:0] add_0_14;
    wire [9-1:0] add_0_15;
    wire [9-1:0] add_0_16;
    wire [9-1:0] add_0_17;
    wire [9-1:0] add_0_18;
    wire [9-1:0] add_0_19;
    wire [9-1:0] add_0_20;
    wire [9-1:0] add_0_21;
    wire [9-1:0] add_0_22;
    wire [9-1:0] add_0_23;
    wire [9-1:0] add_0_24;
    wire [9-1:0] add_0_25;
    wire [9-1:0] add_0_26;
    wire [9-1:0] add_0_27;
    wire [9-1:0] add_0_28;
    wire [9-1:0] add_0_29;
    wire [9-1:0] add_0_30;
    wire [9-1:0] add_0_31;

    wire [10-1:0] add_1_00;
    wire [10-1:0] add_1_01;
    wire [10-1:0] add_1_02;
    wire [10-1:0] add_1_03;
    wire [10-1:0] add_1_04;
    wire [10-1:0] add_1_05;
    wire [10-1:0] add_1_06;
    wire [10-1:0] add_1_07;
    wire [10-1:0] add_1_08;
    wire [10-1:0] add_1_09;
    wire [10-1:0] add_1_10;
    wire [10-1:0] add_1_11;
    wire [10-1:0] add_1_12;
    wire [10-1:0] add_1_13;
    wire [10-1:0] add_1_14;
    wire [10-1:0] add_1_15;

    wire [11-1:0] add_2_0;
    wire [11-1:0] add_2_1;
    wire [11-1:0] add_2_2;
    wire [11-1:0] add_2_3;
    wire [11-1:0] add_2_4;
    wire [11-1:0] add_2_5;
    wire [11-1:0] add_2_6;
    wire [11-1:0] add_2_7;

    wire [12-1:0] add_3_0;
    wire [12-1:0] add_3_1;
    wire [12-1:0] add_3_2;
    wire [12-1:0] add_3_3;

    wire [13-1:0] add_4_0;
    wire [13-1:0] add_4_1;
    //wire [14-1:0] add_5_0 = sad

    assign add_0_00 = ad_00 + ad_01;
    assign add_0_01 = ad_02 + ad_03;
    assign add_0_02 = ad_04 + ad_05;
    assign add_0_03 = ad_06 + ad_07;
    assign add_0_04 = ad_10 + ad_11;
    assign add_0_05 = ad_12 + ad_13;
    assign add_0_06 = ad_14 + ad_15;
    assign add_0_07 = ad_16 + ad_17;
    assign add_0_08 = ad_20 + ad_21;
    assign add_0_09 = ad_22 + ad_23;
    assign add_0_10 = ad_24 + ad_25;
    assign add_0_11 = ad_26 + ad_27;
    assign add_0_12 = ad_30 + ad_31;
    assign add_0_13 = ad_32 + ad_33;
    assign add_0_14 = ad_34 + ad_35;
    assign add_0_15 = ad_36 + ad_37;
    assign add_0_16 = ad_40 + ad_41;
    assign add_0_17 = ad_42 + ad_43;
    assign add_0_18 = ad_44 + ad_45;
    assign add_0_19 = ad_46 + ad_47;
    assign add_0_20 = ad_50 + ad_51;
    assign add_0_21 = ad_52 + ad_53;
    assign add_0_22 = ad_54 + ad_55;
    assign add_0_23 = ad_56 + ad_57;
    assign add_0_24 = ad_60 + ad_61;
    assign add_0_25 = ad_62 + ad_63;
    assign add_0_26 = ad_64 + ad_65;
    assign add_0_27 = ad_66 + ad_67;
    assign add_0_28 = ad_70 + ad_71;
    assign add_0_29 = ad_72 + ad_73;
    assign add_0_30 = ad_74 + ad_75;
    assign add_0_31 = ad_76 + ad_77;

    assign add_1_00 = add_0_00 + add_0_01;
    assign add_1_01 = add_0_02 + add_0_03;
    assign add_1_02 = add_0_04 + add_0_05;
    assign add_1_03 = add_0_06 + add_0_07;
    assign add_1_04 = add_0_08 + add_0_09;
    assign add_1_05 = add_0_10 + add_0_11;
    assign add_1_06 = add_0_12 + add_0_13;
    assign add_1_07 = add_0_14 + add_0_15;
    assign add_1_08 = add_0_16 + add_0_17;
    assign add_1_09 = add_0_18 + add_0_19;
    assign add_1_10 = add_0_20 + add_0_21;
    assign add_1_11 = add_0_22 + add_0_23;
    assign add_1_12 = add_0_24 + add_0_25;
    assign add_1_13 = add_0_26 + add_0_27;
    assign add_1_14 = add_0_28 + add_0_29;
    assign add_1_15 = add_0_30 + add_0_31;

    assign add_2_0 = add_1_00 + add_1_01;
    assign add_2_1 = add_1_02 + add_1_03;
    assign add_2_2 = add_1_04 + add_1_05;
    assign add_2_3 = add_1_06 + add_1_07;
    assign add_2_4 = add_1_08 + add_1_09;
    assign add_2_5 = add_1_10 + add_1_11;
    assign add_2_6 = add_1_12 + add_1_13;
    assign add_2_7 = add_1_14 + add_1_15;

    assign add_3_0 = add_2_0 + add_2_1;
    assign add_3_1 = add_2_2 + add_2_3;
    assign add_3_2 = add_2_4 + add_2_5;
    assign add_3_3 = add_2_6 + add_2_7;

    assign add_4_0 = add_3_0 + add_3_1;
    assign add_4_1 = add_3_2 + add_3_3;

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            sad_data <= 0;
        end
        else begin
            sad_data <= add_4_0 + add_4_1;
        end
    end

endmodule
