module pe (
    input wire [8-1:0] crt_pixel_i,
    input wire [8-1:0] pre_pixel_i,
    output wire [8-1:0] crt_pixel_o,
    output wire [8-1:0] pre_pixel_o,
    output wire [8-1:0] ad 
);
    
endmodule